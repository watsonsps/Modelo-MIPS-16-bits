library ieee;
use ieee.std_logic_1164.all;
use work.all;
use ieee.numeric_std.all;

entity IR is 
	port (
		Write_Reg : in std_logic_vector(15 downto 0);
		Reg_1: out std_logic_vector (15 downto 0)
		);
end IR;

architecture comportamento of IR is

	begin
	process (Write_Reg)
		begin
		case Write_Reg is
		
			-- inicia:
		
			when "0000000000000000" => --0-la-
				Reg_1 <= "0001011100000000";
				
			when "0000000000000001" => --1-addi-
				Reg_1 <= "0001010100000000";
				
			when "0000000000000010" => --2-addi-
				Reg_1 <= "0001011000000000";
				
			when "0000000000000011" => --3-addi-
				Reg_1 <= "0001001000000000";
				
			when "0000000000000100" => --4-addi-
				Reg_1 <= "0001100100000011";
				
			--for1: 
				
			when "0000000000000101" => --5-slti-
				Reg_1 <= "1000000101010011";
				
			when "0000000000000110" => --6-beq
				Reg_1 <= "1001000000000001";
				
			when "0000000000000111" => --7-subi
				Reg_1 <= "1101011001010001";
			
			-- for2:	
				
			when "0000000000001000" => --8-slti
				Reg_1 <= "1000000101100000";
				
			when "0000000000001001" => --9-bne 
				Reg_1 <= "1010010000000001";
				
			when "0000000000001010" => --10-add
				Reg_1 <= "0000100001110110";
				
			when "0000000000001011" => --11-lw 
				Reg_1 <= "0011001110000000";
				
			when "0000000000001100" => --12-lw
				Reg_1 <= "0011010010000001";
				
			when "0000000000001101" => --13-slt
				Reg_1 <= "0111000101000011";
				
			when "0000000000001110" => --14-beq 
				Reg_1 <= "1001100000000001";
				
			-- troca:
				
			when "0000000000001111" => --15-sw
				Reg_1 <= "0100000010000100";
				
			when "0000000000010000" => --16-sw 
				Reg_1 <= "0100000110000011";
				
			-- após a troca: 
				
			when "0000000000010001" => --17-subi
				Reg_1 <= "1101011001100001";
				
			when "0000000000010010" => --18-j 
				Reg_1 <= "1011111111110110";
				
			-- exit2: 
				
			when "0000000000010011" => --19-addi 
				Reg_1 <= "0001010101010001";
				
			when "0000000000010100" => --20-j
				Reg_1 <= "1011111111110001";
				
			when "0000000000010101" => --21-addi
				Reg_1 <= "0001011000000000";
				
			-- exit1: 
				
			when "0000000000010110" => --22-slt 
				Reg_1 <= "0111000101101001";
				
			when "0000000000010111" => --23-beq
				Reg_1 <= "1001110000000001";
				
			when "0000000000011000" => --24-add
				Reg_1 <= "0000100001100111";
				
			when "0000000000011001" => --25-lw 
				Reg_1 <= "0011001110000000";
				
			when "0000000000011010" => --26-add
				Reg_1 <= "0000001000100011";
				
			when "0000000000011011" => --27-addi
				Reg_1 <= "0001011001100001";
				
			when "0000000000011100" => --28-j
				Reg_1 <= "1011111111111010";
				
			
			when "0000000000011101" => --29-sw
				Reg_1 <= "0100001101110010";
				--exit_loop_pre:
				
			when "0000000000011110" => --30-regIN-lw
				Reg_1 <= "0011000101111110";
				
			when "0000000000011111" => --30-regIN-lw
				Reg_1 <= "0011001000010000";
				
			when "0000000000100000" => --31-regOUT-sw
				Reg_1 <= "0100111101110010";
				
			-- exit_loop:
			when others => --34-loop para debug final
				Reg_1 <= "1011111111111101";
					
		end case;	
	end process;
end comportamento;